module fa_ha(a,b,c,sum,carry);
input a,b,c;
output sum,carry;



endmodule
