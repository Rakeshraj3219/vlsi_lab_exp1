module hs(a,b,difference,borrow);
input a,b;
output difference,borrow;



endmodule
